package ahb_vga_font_map;

	string font_map [128] = {
		" ",
		"☺",
		"☻",
		"♥",
		"◆",
		"♣",
		"♠",
		"·",
		" ",
		"○",
		" ",
		"♂",
		"♀",
		" ",
		"♬",
		"☼",
		"⏵",
		"⏴",
		"↕",
		"‼",
		"¶",
		"§",
		"⏹",
		"↨",
		"↑",
		"↓",
		"→",
		"←",
		"∟",
		"↔",
		"▲",
		"▼",
		" ",
		"❢",
		"\"",
		"#",
		"$",
		"%",
		"&",
		"'",
		"(",
		")",
		"*",
		"+",
		",",
		"-",
		".",
		"/",
		"0",
		"1",
		"2",
		"3",
		"4",
		"5",
		"6",
		"7",
		"8",
		"9",
		":",
		";",
		"<",
		"=",
		">",
		"?",
		"@",
		"A",
		"B",
		"C",
		"D",
		"E",
		"F",
		"G",
		"H",
		"I",
		"J",
		"K",
		"L",
		"M",
		"N",
		"O",
		"P",
		"Q",
		"R",
		"S",
		"T",
		"U",
		"V",
		"W",
		"X",
		"Y",
		"Z",
		"[",
		"\\",
		"]",
		"^",
		"_",
		"`",
		"a",
		"b",
		"c",
		"d",
		"e",
		"f",
		"g",
		"h",
		"i",
		"j",
		"k",
		"l",
		"m",
		"n",
		"o",
		"p",
		"q",
		"r",
		"s",
		"t",
		"u",
		"v",
		"w",
		"x",
		"y",
		"z",
		"{",
		"|",
		"}",
		"~",
		"🏠"
	};


  function int font_lookup(logic [10:0] addr);
    case (addr)
         //code x00
         11'h000: return 8'b00000000; //
         11'h001: return 8'b00000000; //
         11'h002: return 8'b00000000; //
         11'h003: return 8'b00000000; //
         11'h004: return 8'b00000000; //
         11'h005: return 8'b00000000; //
         11'h006: return 8'b00000000; //
         11'h007: return 8'b00000000; //
         11'h008: return 8'b00000000; //
         11'h009: return 8'b00000000; //
         11'h00a: return 8'b00000000; //
         11'h00b: return 8'b00000000; //
         11'h00c: return 8'b00000000; //
         11'h00d: return 8'b00000000; //
         11'h00e: return 8'b00000000; //
         11'h00f: return 8'b00000000; //
         //code x01
         11'h010: return 8'b00000000; //
         11'h011: return 8'b00000000; //
         11'h012: return 8'b01111110; //  ******
         11'h013: return 8'b10000001; // *      *
         11'h014: return 8'b10100101; // * *  * *
         11'h015: return 8'b10000001; // *      *
         11'h016: return 8'b10000001; // *      *
         11'h017: return 8'b10111101; // * **** *
         11'h018: return 8'b10011001; // *  **  *
         11'h019: return 8'b10000001; // *      *
         11'h01a: return 8'b10000001; // *      *
         11'h01b: return 8'b01111110; //  ******
         11'h01c: return 8'b00000000; //
         11'h01d: return 8'b00000000; //
         11'h01e: return 8'b00000000; //
         11'h01f: return 8'b00000000; //
         //code x02
         11'h020: return 8'b00000000; //
         11'h021: return 8'b00000000; //
         11'h022: return 8'b01111110; //  ******
         11'h023: return 8'b11111111; // ********
         11'h024: return 8'b11011011; // ** ** **
         11'h025: return 8'b11111111; // ********
         11'h026: return 8'b11111111; // ********
         11'h027: return 8'b11000011; // **    **
         11'h028: return 8'b11100111; // ***  ***
         11'h029: return 8'b11111111; // ********
         11'h02a: return 8'b11111111; // ********
         11'h02b: return 8'b01111110; //  ******
         11'h02c: return 8'b00000000; //
         11'h02d: return 8'b00000000; //
         11'h02e: return 8'b00000000; //
         11'h02f: return 8'b00000000; //
         //code x03
         11'h030: return 8'b00000000; //
         11'h031: return 8'b00000000; //
         11'h032: return 8'b00000000; //
         11'h033: return 8'b00000000; //
         11'h034: return 8'b01101100; //  ** **
         11'h035: return 8'b11111110; // *******
         11'h036: return 8'b11111110; // *******
         11'h037: return 8'b11111110; // *******
         11'h038: return 8'b11111110; // *******
         11'h039: return 8'b01111100; //  *****
         11'h03a: return 8'b00111000; //   ***
         11'h03b: return 8'b00010000; //    *
         11'h03c: return 8'b00000000; //
         11'h03d: return 8'b00000000; //
         11'h03e: return 8'b00000000; //
         11'h03f: return 8'b00000000; //
         //code x04
         11'h040: return 8'b00000000; //
         11'h041: return 8'b00000000; //
         11'h042: return 8'b00000000; //
         11'h043: return 8'b00000000; //
         11'h044: return 8'b00010000; //    *
         11'h045: return 8'b00111000; //   ***
         11'h046: return 8'b01111100; //  *****
         11'h047: return 8'b11111110; // *******
         11'h048: return 8'b01111100; //  *****
         11'h049: return 8'b00111000; //   ***
         11'h04a: return 8'b00010000; //    *
         11'h04b: return 8'b00000000; //
         11'h04c: return 8'b00000000; //
         11'h04d: return 8'b00000000; //
         11'h04e: return 8'b00000000; //
         11'h04f: return 8'b00000000; //
         //code x05
         11'h050: return 8'b00000000; //
         11'h051: return 8'b00000000; //
         11'h052: return 8'b00000000; //
         11'h053: return 8'b00011000; //    **
         11'h054: return 8'b00111100; //   ****
         11'h055: return 8'b00111100; //   ****
         11'h056: return 8'b11100111; // ***  ***
         11'h057: return 8'b11100111; // ***  ***
         11'h058: return 8'b11100111; // ***  ***
         11'h059: return 8'b00011000; //    **
         11'h05a: return 8'b00011000; //    **
         11'h05b: return 8'b00111100; //   ****
         11'h05c: return 8'b00000000; //
         11'h05d: return 8'b00000000; //
         11'h05e: return 8'b00000000; //
         11'h05f: return 8'b00000000; //
         //code x06
         11'h060: return 8'b00000000; //
         11'h061: return 8'b00000000; //
         11'h062: return 8'b00000000; //
         11'h063: return 8'b00011000; //    **
         11'h064: return 8'b00111100; //   ****
         11'h065: return 8'b01111110; //  ******
         11'h066: return 8'b11111111; // ********
         11'h067: return 8'b11111111; // ********
         11'h068: return 8'b01111110; //  ******
         11'h069: return 8'b00011000; //    **
         11'h06a: return 8'b00011000; //    **
         11'h06b: return 8'b00111100; //   ****
         11'h06c: return 8'b00000000; //
         11'h06d: return 8'b00000000; //
         11'h06e: return 8'b00000000; //
         11'h06f: return 8'b00000000; //
         //code x07
         11'h070: return 8'b00000000; //
         11'h071: return 8'b00000000; //
         11'h072: return 8'b00000000; //
         11'h073: return 8'b00000000; //
         11'h074: return 8'b00000000; //
         11'h075: return 8'b00000000; //
         11'h076: return 8'b00011000; //    **
         11'h077: return 8'b00111100; //   ****
         11'h078: return 8'b00111100; //   ****
         11'h079: return 8'b00011000; //    **
         11'h07a: return 8'b00000000; //
         11'h07b: return 8'b00000000; //
         11'h07c: return 8'b00000000; //
         11'h07d: return 8'b00000000; //
         11'h07e: return 8'b00000000; //
         11'h07f: return 8'b00000000; //
         //code x08
         11'h080: return 8'b00000000; //
         11'h081: return 8'b00000000; //
         11'h082: return 8'b00000000; //
         11'h083: return 8'b00000000; //
         11'h084: return 8'b00000000; //
         11'h085: return 8'b00000000; //
         11'h086: return 8'b00000000; //
         11'h087: return 8'b00000000; //
         11'h088: return 8'b00000000; //
         11'h089: return 8'b00000000; //
         11'h08a: return 8'b00000000; //
         11'h08b: return 8'b00000000; //
         11'h08c: return 8'b00000000; //
         11'h08d: return 8'b00000000; //
         11'h08e: return 8'b00000000; //
         11'h08f: return 8'b00000000; //
         //code x09
         11'h090: return 8'b00000000; //
         11'h091: return 8'b00000000; //
         11'h092: return 8'b00000000; //
         11'h093: return 8'b00000000; //
         11'h094: return 8'b00000000; //
         11'h095: return 8'b00111100; //   ****
         11'h096: return 8'b01100110; //  **  **
         11'h097: return 8'b01000010; //  *    *
         11'h098: return 8'b01000010; //  *    *
         11'h099: return 8'b01100110; //  **  **
         11'h09a: return 8'b00111100; //   ****
         11'h09b: return 8'b00000000; //
         11'h09c: return 8'b00000000; //
         11'h09d: return 8'b00000000; //
         11'h09e: return 8'b00000000; //
         11'h09f: return 8'b00000000; //
         //code x0a
         11'h0a0: return 8'b00000000; //
         11'h0a1: return 8'b00000000; //
         11'h0a2: return 8'b00000000; //
         11'h0a3: return 8'b00000000; //
         11'h0a4: return 8'b00000000; //
         11'h0a5: return 8'b00000000; //
         11'h0a6: return 8'b00000000; //
         11'h0a7: return 8'b00000000; //
         11'h0a8: return 8'b00000000; //
         11'h0a9: return 8'b00000000; //
         11'h0aa: return 8'b00000000; //
         11'h0ab: return 8'b00000000; //
         11'h0ac: return 8'b00000000; //
         11'h0ad: return 8'b00000000; //
         11'h0ae: return 8'b00000000; //
         11'h0af: return 8'b00000000; //
         //code x0b
         11'h0b0: return 8'b00000000; //
         11'h0b1: return 8'b00000000; //
         11'h0b2: return 8'b00011110; //    ****
         11'h0b3: return 8'b00001110; //     ***
         11'h0b4: return 8'b00011010; //    ** *
         11'h0b5: return 8'b00110010; //   **  *
         11'h0b6: return 8'b01111000; //  ****
         11'h0b7: return 8'b11001100; // **  **
         11'h0b8: return 8'b11001100; // **  **
         11'h0b9: return 8'b11001100; // **  **
         11'h0ba: return 8'b11001100; // **  **
         11'h0bb: return 8'b01111000; //  ****
         11'h0bc: return 8'b00000000; //
         11'h0bd: return 8'b00000000; //
         11'h0be: return 8'b00000000; //
         11'h0bf: return 8'b00000000; //
         //code x0c
         11'h0c0: return 8'b00000000; //
         11'h0c1: return 8'b00000000; //
         11'h0c2: return 8'b00111100; //   ****
         11'h0c3: return 8'b01100110; //  **  **
         11'h0c4: return 8'b01100110; //  **  **
         11'h0c5: return 8'b01100110; //  **  **
         11'h0c6: return 8'b01100110; //  **  **
         11'h0c7: return 8'b00111100; //   ****
         11'h0c8: return 8'b00011000; //    **
         11'h0c9: return 8'b01111110; //  ******
         11'h0ca: return 8'b00011000; //    **
         11'h0cb: return 8'b00011000; //    **
         11'h0cc: return 8'b00000000; //
         11'h0cd: return 8'b00000000; //
         11'h0ce: return 8'b00000000; //
         11'h0cf: return 8'b00000000; //
         //code x0d
         11'h0d0: return 8'b00000000; //
         11'h0d1: return 8'b00000000; //
         11'h0d2: return 8'b00000000; //
         11'h0d3: return 8'b00000000; //
         11'h0d4: return 8'b00000000; //
         11'h0d5: return 8'b00000000; //
         11'h0d6: return 8'b00000000; //
         11'h0d7: return 8'b00000000; //
         11'h0d8: return 8'b00000000; //
         11'h0d9: return 8'b00000000; //
         11'h0da: return 8'b00000000; //
         11'h0db: return 8'b00000000; //
         11'h0dc: return 8'b00000000; //
         11'h0dd: return 8'b00000000; //
         11'h0de: return 8'b00000000; //
         11'h0df: return 8'b00000000; //
         //code x0e
         11'h0e0: return 8'b00000000; //
         11'h0e1: return 8'b00000000; //
         11'h0e2: return 8'b01111111; //  *******
         11'h0e3: return 8'b01100011; //  **   **
         11'h0e4: return 8'b01111111; //  *******
         11'h0e5: return 8'b01100011; //  **   **
         11'h0e6: return 8'b01100011; //  **   **
         11'h0e7: return 8'b01100011; //  **   **
         11'h0e8: return 8'b01100011; //  **   **
         11'h0e9: return 8'b01100111; //  **  ***
         11'h0ea: return 8'b11100111; // ***  ***
         11'h0eb: return 8'b11100110; // ***  **
         11'h0ec: return 8'b11000000; // **
         11'h0ed: return 8'b00000000; //
         11'h0ee: return 8'b00000000; //
         11'h0ef: return 8'b00000000; //
         //code x0f
         11'h0f0: return 8'b00000000; //
         11'h0f1: return 8'b00000000; //
         11'h0f2: return 8'b00000000; //
         11'h0f3: return 8'b00011000; //    **
         11'h0f4: return 8'b00011000; //    **
         11'h0f5: return 8'b11011011; // ** ** **
         11'h0f6: return 8'b00111100; //   ****
         11'h0f7: return 8'b11100111; // ***  ***
         11'h0f8: return 8'b00111100; //   ****
         11'h0f9: return 8'b11011011; // ** ** **
         11'h0fa: return 8'b00011000; //    **
         11'h0fb: return 8'b00011000; //    **
         11'h0fc: return 8'b00000000; //
         11'h0fd: return 8'b00000000; //
         11'h0fe: return 8'b00000000; //
         11'h0ff: return 8'b00000000; //
         //code x10
         11'h100: return 8'b00000000; //
         11'h101: return 8'b10000000; // *
         11'h102: return 8'b11000000; // **
         11'h103: return 8'b11100000; // ***
         11'h104: return 8'b11110000; // ****
         11'h105: return 8'b11111000; // *****
         11'h106: return 8'b11111110; // *******
         11'h107: return 8'b11111000; // *****
         11'h108: return 8'b11110000; // ****
         11'h109: return 8'b11100000; // ***
         11'h10a: return 8'b11000000; // **
         11'h10b: return 8'b10000000; // *
         11'h10c: return 8'b00000000; //
         11'h10d: return 8'b00000000; //
         11'h10e: return 8'b00000000; //
         11'h10f: return 8'b00000000; //
         //code x11
         11'h110: return 8'b00000000; //
         11'h111: return 8'b00000010; //       *
         11'h112: return 8'b00000110; //      **
         11'h113: return 8'b00001110; //     ***
         11'h114: return 8'b00011110; //    ****
         11'h115: return 8'b00111110; //   *****
         11'h116: return 8'b11111110; // *******
         11'h117: return 8'b00111110; //   *****
         11'h118: return 8'b00011110; //    ****
         11'h119: return 8'b00001110; //     ***
         11'h11a: return 8'b00000110; //      **
         11'h11b: return 8'b00000010; //       *
         11'h11c: return 8'b00000000; //
         11'h11d: return 8'b00000000; //
         11'h11e: return 8'b00000000; //
         11'h11f: return 8'b00000000; //
         //code x12
         11'h120: return 8'b00000000; //
         11'h121: return 8'b00000000; //
         11'h122: return 8'b00011000; //    **
         11'h123: return 8'b00111100; //   ****
         11'h124: return 8'b01111110; //  ******
         11'h125: return 8'b00011000; //    **
         11'h126: return 8'b00011000; //    **
         11'h127: return 8'b00011000; //    **
         11'h128: return 8'b01111110; //  ******
         11'h129: return 8'b00111100; //   ****
         11'h12a: return 8'b00011000; //    **
         11'h12b: return 8'b00000000; //
         11'h12c: return 8'b00000000; //
         11'h12d: return 8'b00000000; //
         11'h12e: return 8'b00000000; //
         11'h12f: return 8'b00000000; //
         //code x13
         11'h130: return 8'b00000000; //
         11'h131: return 8'b00000000; //
         11'h132: return 8'b01100110; //  **  **
         11'h133: return 8'b01100110; //  **  **
         11'h134: return 8'b01100110; //  **  **
         11'h135: return 8'b01100110; //  **  **
         11'h136: return 8'b01100110; //  **  **
         11'h137: return 8'b01100110; //  **  **
         11'h138: return 8'b01100110; //  **  **
         11'h139: return 8'b00000000; //
         11'h13a: return 8'b01100110; //  **  **
         11'h13b: return 8'b01100110; //  **  **
         11'h13c: return 8'b00000000; //
         11'h13d: return 8'b00000000; //
         11'h13e: return 8'b00000000; //
         11'h13f: return 8'b00000000; //
         //code x14
         11'h140: return 8'b00000000; //
         11'h141: return 8'b00000000; //
         11'h142: return 8'b01111111; //  *******
         11'h143: return 8'b11011011; // ** ** **
         11'h144: return 8'b11011011; // ** ** **
         11'h145: return 8'b11011011; // ** ** **
         11'h146: return 8'b01111011; //  **** **
         11'h147: return 8'b00011011; //    ** **
         11'h148: return 8'b00011011; //    ** **
         11'h149: return 8'b00011011; //    ** **
         11'h14a: return 8'b00011011; //    ** **
         11'h14b: return 8'b00011011; //    ** **
         11'h14c: return 8'b00000000; //
         11'h14d: return 8'b00000000; //
         11'h14e: return 8'b00000000; //
         11'h14f: return 8'b00000000; //
         //code x15
         11'h150: return 8'b00000000; //
         11'h151: return 8'b01111100; //  *****
         11'h152: return 8'b11000110; // **   **
         11'h153: return 8'b01100000; //  **
         11'h154: return 8'b00111000; //   ***
         11'h155: return 8'b01101100; //  ** **
         11'h156: return 8'b11000110; // **   **
         11'h157: return 8'b11000110; // **   **
         11'h158: return 8'b01101100; //  ** **
         11'h159: return 8'b00111000; //   ***
         11'h15a: return 8'b00001100; //     **
         11'h15b: return 8'b11000110; // **   **
         11'h15c: return 8'b01111100; //  *****
         11'h15d: return 8'b00000000; //
         11'h15e: return 8'b00000000; //
         11'h15f: return 8'b00000000; //
         //code x16
         11'h160: return 8'b00000000; //
         11'h161: return 8'b00000000; //
         11'h162: return 8'b00000000; //
         11'h163: return 8'b00000000; //
         11'h164: return 8'b00000000; //
         11'h165: return 8'b00000000; //
         11'h166: return 8'b00000000; //
         11'h167: return 8'b00000000; //
         11'h168: return 8'b11111110; // *******
         11'h169: return 8'b11111110; // *******
         11'h16a: return 8'b11111110; // *******
         11'h16b: return 8'b11111110; // *******
         11'h16c: return 8'b00000000; //
         11'h16d: return 8'b00000000; //
         11'h16e: return 8'b00000000; //
         11'h16f: return 8'b00000000; //
         //code x17
         11'h170: return 8'b00000000; //
         11'h171: return 8'b00000000; //
         11'h172: return 8'b00011000; //    **
         11'h173: return 8'b00111100; //   ****
         11'h174: return 8'b01111110; //  ******
         11'h175: return 8'b00011000; //    **
         11'h176: return 8'b00011000; //    **
         11'h177: return 8'b00011000; //    **
         11'h178: return 8'b01111110; //  ******
         11'h179: return 8'b00111100; //   ****
         11'h17a: return 8'b00011000; //    **
         11'h17b: return 8'b01111110; //  ******
         11'h17c: return 8'b00110000; //
         11'h17d: return 8'b00000000; //
         11'h17e: return 8'b00000000; //
         11'h17f: return 8'b00000000; //
         //code x18
         11'h180: return 8'b00000000; //
         11'h181: return 8'b00000000; //
         11'h182: return 8'b00011000; //    **
         11'h183: return 8'b00111100; //   ****
         11'h184: return 8'b01111110; //  ******
         11'h185: return 8'b00011000; //    **
         11'h186: return 8'b00011000; //    **
         11'h187: return 8'b00011000; //    **
         11'h188: return 8'b00011000; //    **
         11'h189: return 8'b00011000; //    **
         11'h18a: return 8'b00011000; //    **
         11'h18b: return 8'b00011000; //    **
         11'h18c: return 8'b00000000; //
         11'h18d: return 8'b00000000; //
         11'h18e: return 8'b00000000; //
         11'h18f: return 8'b00000000; //
         //code x19
         11'h190: return 8'b00000000; //
         11'h191: return 8'b00000000; //
         11'h192: return 8'b00011000; //    **
         11'h193: return 8'b00011000; //    **
         11'h194: return 8'b00011000; //    **
         11'h195: return 8'b00011000; //    **
         11'h196: return 8'b00011000; //    **
         11'h197: return 8'b00011000; //    **
         11'h198: return 8'b00011000; //    **
         11'h199: return 8'b01111110; //  ******
         11'h19a: return 8'b00111100; //   ****
         11'h19b: return 8'b00011000; //    **
         11'h19c: return 8'b00000000; //
         11'h19d: return 8'b00000000; //
         11'h19e: return 8'b00000000; //
         11'h19f: return 8'b00000000; //
         //code x1a
         11'h1a0: return 8'b00000000; //
         11'h1a1: return 8'b00000000; //
         11'h1a2: return 8'b00000000; //
         11'h1a3: return 8'b00000000; //
         11'h1a4: return 8'b00000000; //
         11'h1a5: return 8'b00011000; //    **
         11'h1a6: return 8'b00001100; //     **
         11'h1a7: return 8'b11111110; // *******
         11'h1a8: return 8'b00001100; //     **
         11'h1a9: return 8'b00011000; //    **
         11'h1aa: return 8'b00000000; //
         11'h1ab: return 8'b00000000; //
         11'h1ac: return 8'b00000000; //
         11'h1ad: return 8'b00000000; //
         11'h1ae: return 8'b00000000; //
         11'h1af: return 8'b00000000; //
         //code x1b
         11'h1b0: return 8'b00000000; //
         11'h1b1: return 8'b00000000; //
         11'h1b2: return 8'b00000000; //
         11'h1b3: return 8'b00000000; //
         11'h1b4: return 8'b00000000; //
         11'h1b5: return 8'b00110000; //   **
         11'h1b6: return 8'b01100000; //  **
         11'h1b7: return 8'b11111110; // *******
         11'h1b8: return 8'b01100000; //  **
         11'h1b9: return 8'b00110000; //   **
         11'h1ba: return 8'b00000000; //
         11'h1bb: return 8'b00000000; //
         11'h1bc: return 8'b00000000; //
         11'h1bd: return 8'b00000000; //
         11'h1be: return 8'b00000000; //
         11'h1bf: return 8'b00000000; //
         //code x1c
         11'h1c0: return 8'b00000000; //
         11'h1c1: return 8'b00000000; //
         11'h1c2: return 8'b00000000; //
         11'h1c3: return 8'b00000000; //
         11'h1c4: return 8'b00000000; //
         11'h1c5: return 8'b00000000; //
         11'h1c6: return 8'b11000000; // **
         11'h1c7: return 8'b11000000; // **
         11'h1c8: return 8'b11000000; // **
         11'h1c9: return 8'b11111110; // *******
         11'h1ca: return 8'b00000000; //
         11'h1cb: return 8'b00000000; //
         11'h1cc: return 8'b00000000; //
         11'h1cd: return 8'b00000000; //
         11'h1ce: return 8'b00000000; //
         11'h1cf: return 8'b00000000; //
         //code x1d
         11'h1d0: return 8'b00000000; //
         11'h1d1: return 8'b00000000; //
         11'h1d2: return 8'b00000000; //
         11'h1d3: return 8'b00000000; //
         11'h1d4: return 8'b00000000; //
         11'h1d5: return 8'b00100100; //   *  *
         11'h1d6: return 8'b01100110; //  **  **
         11'h1d7: return 8'b11111111; // ********
         11'h1d8: return 8'b01100110; //  **  **
         11'h1d9: return 8'b00100100; //   *  *
         11'h1da: return 8'b00000000; //
         11'h1db: return 8'b00000000; //
         11'h1dc: return 8'b00000000; //
         11'h1dd: return 8'b00000000; //
         11'h1de: return 8'b00000000; //
         11'h1df: return 8'b00000000; //
         //code x1e
         11'h1e0: return 8'b00000000; //
         11'h1e1: return 8'b00000000; //
         11'h1e2: return 8'b00000000; //
         11'h1e3: return 8'b00000000; //
         11'h1e4: return 8'b00010000; //    *
         11'h1e5: return 8'b00111000; //   ***
         11'h1e6: return 8'b00111000; //   ***
         11'h1e7: return 8'b01111100; //  *****
         11'h1e8: return 8'b01111100; //  *****
         11'h1e9: return 8'b11111110; // *******
         11'h1ea: return 8'b11111110; // *******
         11'h1eb: return 8'b00000000; //
         11'h1ec: return 8'b00000000; //
         11'h1ed: return 8'b00000000; //
         11'h1ee: return 8'b00000000; //
         11'h1ef: return 8'b00000000; //
         //code x1f
         11'h1f0: return 8'b00000000; //
         11'h1f1: return 8'b00000000; //
         11'h1f2: return 8'b00000000; //
         11'h1f3: return 8'b00000000; //
         11'h1f4: return 8'b11111110; // *******
         11'h1f5: return 8'b11111110; // *******
         11'h1f6: return 8'b01111100; //  *****
         11'h1f7: return 8'b01111100; //  *****
         11'h1f8: return 8'b00111000; //   ***
         11'h1f9: return 8'b00111000; //   ***
         11'h1fa: return 8'b00010000; //    *
         11'h1fb: return 8'b00000000; //
         11'h1fc: return 8'b00000000; //
         11'h1fd: return 8'b00000000; //
         11'h1fe: return 8'b00000000; //
         11'h1ff: return 8'b00000000; //
         //code x20
         11'h200: return 8'b00000000; //
         11'h201: return 8'b00000000; //
         11'h202: return 8'b00000000; //
         11'h203: return 8'b00000000; //
         11'h204: return 8'b00000000; //
         11'h205: return 8'b00000000; //
         11'h206: return 8'b00000000; //
         11'h207: return 8'b00000000; //
         11'h208: return 8'b00000000; //
         11'h209: return 8'b00000000; //
         11'h20a: return 8'b00000000; //
         11'h20b: return 8'b00000000; //
         11'h20c: return 8'b00000000; //
         11'h20d: return 8'b00000000; //
         11'h20e: return 8'b00000000; //
         11'h20f: return 8'b00000000; //
         //code x21
         11'h210: return 8'b00000000; //
         11'h211: return 8'b00000000; //
         11'h212: return 8'b00011000; //    **
         11'h213: return 8'b00111100; //   ****
         11'h214: return 8'b00111100; //   ****
         11'h215: return 8'b00111100; //   ****
         11'h216: return 8'b00011000; //    **
         11'h217: return 8'b00011000; //    **
         11'h218: return 8'b00011000; //    **
         11'h219: return 8'b00000000; //
         11'h21a: return 8'b00011000; //    **
         11'h21b: return 8'b00011000; //    **
         11'h21c: return 8'b00000000; //
         11'h21d: return 8'b00000000; //
         11'h21e: return 8'b00000000; //
         11'h21f: return 8'b00000000; //
         //code x22
         11'h220: return 8'b00000000; //
         11'h221: return 8'b01100110; //  **  **
         11'h222: return 8'b01100110; //  **  **
         11'h223: return 8'b01100110; //  **  **
         11'h224: return 8'b00100100; //   *  *
         11'h225: return 8'b00000000; //
         11'h226: return 8'b00000000; //
         11'h227: return 8'b00000000; //
         11'h228: return 8'b00000000; //
         11'h229: return 8'b00000000; //
         11'h22a: return 8'b00000000; //
         11'h22b: return 8'b00000000; //
         11'h22c: return 8'b00000000; //
         11'h22d: return 8'b00000000; //
         11'h22e: return 8'b00000000; //
         11'h22f: return 8'b00000000; //
         //code x23
         11'h230: return 8'b00000000; //
         11'h231: return 8'b00000000; //
         11'h232: return 8'b00000000; //
         11'h233: return 8'b01101100; //  ** **
         11'h234: return 8'b01101100; //  ** **
         11'h235: return 8'b11111110; // *******
         11'h236: return 8'b01101100; //  ** **
         11'h237: return 8'b01101100; //  ** **
         11'h238: return 8'b01101100; //  ** **
         11'h239: return 8'b11111110; // *******
         11'h23a: return 8'b01101100; //  ** **
         11'h23b: return 8'b01101100; //  ** **
         11'h23c: return 8'b00000000; //
         11'h23d: return 8'b00000000; //
         11'h23e: return 8'b00000000; //
         11'h23f: return 8'b00000000; //
         //code x24
         11'h240: return 8'b00011000; //     **
         11'h241: return 8'b00011000; //     **
         11'h242: return 8'b01111100; //   *****
         11'h243: return 8'b11000110; //  **   **
         11'h244: return 8'b11000010; //  **    *
         11'h245: return 8'b11000000; //  **
         11'h246: return 8'b01111100; //   *****
         11'h247: return 8'b00000110; //       **
         11'h248: return 8'b00000110; //       **
         11'h249: return 8'b10000110; //  *    **
         11'h24a: return 8'b11000110; //  **   **
         11'h24b: return 8'b01111100; //   *****
         11'h24c: return 8'b00011000; //     **
         11'h24d: return 8'b00011000; //     **
         11'h24e: return 8'b00000000; //
         11'h24f: return 8'b00000000; //
         //code x25
         11'h250: return 8'b00000000; //
         11'h251: return 8'b00000000; //
         11'h252: return 8'b00000000; //
         11'h253: return 8'b00000000; //
         11'h254: return 8'b11000010; // **    *
         11'h255: return 8'b11000110; // **   **
         11'h256: return 8'b00001100; //     **
         11'h257: return 8'b00011000; //    **
         11'h258: return 8'b00110000; //   **
         11'h259: return 8'b01100000; //  **
         11'h25a: return 8'b11000110; // **   **
         11'h25b: return 8'b10000110; // *    **
         11'h25c: return 8'b00000000; //
         11'h25d: return 8'b00000000; //
         11'h25e: return 8'b00000000; //
         11'h25f: return 8'b00000000; //
         //code x26
         11'h260: return 8'b00000000; //
         11'h261: return 8'b00000000; //
         11'h262: return 8'b00111000; //   ***
         11'h263: return 8'b01101100; //  ** **
         11'h264: return 8'b01101100; //  ** **
         11'h265: return 8'b00111000; //   ***
         11'h266: return 8'b01110110; //  *** **
         11'h267: return 8'b11011100; // ** ***
         11'h268: return 8'b11001100; // **  **
         11'h269: return 8'b11001100; // **  **
         11'h26a: return 8'b11001100; // **  **
         11'h26b: return 8'b01110110; //  *** **
         11'h26c: return 8'b00000000; //
         11'h26d: return 8'b00000000; //
         11'h26e: return 8'b00000000; //
         11'h26f: return 8'b00000000; //
         //code x27
         11'h270: return 8'b00000000; //
         11'h271: return 8'b00110000; //   **
         11'h272: return 8'b00110000; //   **
         11'h273: return 8'b00110000; //   **
         11'h274: return 8'b01100000; //  **
         11'h275: return 8'b00000000; //
         11'h276: return 8'b00000000; //
         11'h277: return 8'b00000000; //
         11'h278: return 8'b00000000; //
         11'h279: return 8'b00000000; //
         11'h27a: return 8'b00000000; //
         11'h27b: return 8'b00000000; //
         11'h27c: return 8'b00000000; //
         11'h27d: return 8'b00000000; //
         11'h27e: return 8'b00000000; //
         11'h27f: return 8'b00000000; //
         //code x28
         11'h280: return 8'b00000000; //
         11'h281: return 8'b00000000; //
         11'h282: return 8'b00001100; //     **
         11'h283: return 8'b00011000; //    **
         11'h284: return 8'b00110000; //   **
         11'h285: return 8'b00110000; //   **
         11'h286: return 8'b00110000; //   **
         11'h287: return 8'b00110000; //   **
         11'h288: return 8'b00110000; //   **
         11'h289: return 8'b00110000; //   **
         11'h28a: return 8'b00011000; //    **
         11'h28b: return 8'b00001100; //     **
         11'h28c: return 8'b00000000; //
         11'h28d: return 8'b00000000; //
         11'h28e: return 8'b00000000; //
         11'h28f: return 8'b00000000; //
         //code x29
         11'h290: return 8'b00000000; //
         11'h291: return 8'b00000000; //
         11'h292: return 8'b00110000; //   **
         11'h293: return 8'b00011000; //    **
         11'h294: return 8'b00001100; //     **
         11'h295: return 8'b00001100; //     **
         11'h296: return 8'b00001100; //     **
         11'h297: return 8'b00001100; //     **
         11'h298: return 8'b00001100; //     **
         11'h299: return 8'b00001100; //     **
         11'h29a: return 8'b00011000; //    **
         11'h29b: return 8'b00110000; //   **
         11'h29c: return 8'b00000000; //
         11'h29d: return 8'b00000000; //
         11'h29e: return 8'b00000000; //
         11'h29f: return 8'b00000000; //
         //code x2a
         11'h2a0: return 8'b00000000; //
         11'h2a1: return 8'b00000000; //
         11'h2a2: return 8'b00000000; //
         11'h2a3: return 8'b00000000; //
         11'h2a4: return 8'b00000000; //
         11'h2a5: return 8'b01100110; //  **  **
         11'h2a6: return 8'b00111100; //   ****
         11'h2a7: return 8'b11111111; // ********
         11'h2a8: return 8'b00111100; //   ****
         11'h2a9: return 8'b01100110; //  **  **
         11'h2aa: return 8'b00000000; //
         11'h2ab: return 8'b00000000; //
         11'h2ac: return 8'b00000000; //
         11'h2ad: return 8'b00000000; //
         11'h2ae: return 8'b00000000; //
         11'h2af: return 8'b00000000; //
         //code x2b
         11'h2b0: return 8'b00000000; //
         11'h2b1: return 8'b00000000; //
         11'h2b2: return 8'b00000000; //
         11'h2b3: return 8'b00000000; //
         11'h2b4: return 8'b00000000; //
         11'h2b5: return 8'b00011000; //    **
         11'h2b6: return 8'b00011000; //    **
         11'h2b7: return 8'b01111110; //  ******
         11'h2b8: return 8'b00011000; //    **
         11'h2b9: return 8'b00011000; //    **
         11'h2ba: return 8'b00000000; //
         11'h2bb: return 8'b00000000; //
         11'h2bc: return 8'b00000000; //
         11'h2bd: return 8'b00000000; //
         11'h2be: return 8'b00000000; //
         11'h2bf: return 8'b00000000; //
         //code x2c
         11'h2c0: return 8'b00000000; //
         11'h2c1: return 8'b00000000; //
         11'h2c2: return 8'b00000000; //
         11'h2c3: return 8'b00000000; //
         11'h2c4: return 8'b00000000; //
         11'h2c5: return 8'b00000000; //
         11'h2c6: return 8'b00000000; //
         11'h2c7: return 8'b00000000; //
         11'h2c8: return 8'b00000000; //
         11'h2c9: return 8'b00011000; //    **
         11'h2ca: return 8'b00011000; //    **
         11'h2cb: return 8'b00011000; //    **
         11'h2cc: return 8'b00110000; //   **
         11'h2cd: return 8'b00000000; //
         11'h2ce: return 8'b00000000; //
         11'h2cf: return 8'b00000000; //
         //code x2d
         11'h2d0: return 8'b00000000; //
         11'h2d1: return 8'b00000000; //
         11'h2d2: return 8'b00000000; //
         11'h2d3: return 8'b00000000; //
         11'h2d4: return 8'b00000000; //
         11'h2d5: return 8'b00000000; //
         11'h2d6: return 8'b00000000; //
         11'h2d7: return 8'b01111110; //  ******
         11'h2d8: return 8'b00000000; //
         11'h2d9: return 8'b00000000; //
         11'h2da: return 8'b00000000; //
         11'h2db: return 8'b00000000; //
         11'h2dc: return 8'b00000000; //
         11'h2dd: return 8'b00000000; //
         11'h2de: return 8'b00000000; //
         11'h2df: return 8'b00000000; //
         //code x2e
         11'h2e0: return 8'b00000000; //
         11'h2e1: return 8'b00000000; //
         11'h2e2: return 8'b00000000; //
         11'h2e3: return 8'b00000000; //
         11'h2e4: return 8'b00000000; //
         11'h2e5: return 8'b00000000; //
         11'h2e6: return 8'b00000000; //
         11'h2e7: return 8'b00000000; //
         11'h2e8: return 8'b00000000; //
         11'h2e9: return 8'b00000000; //
         11'h2ea: return 8'b00011000; //    **
         11'h2eb: return 8'b00011000; //    **
         11'h2ec: return 8'b00000000; //
         11'h2ed: return 8'b00000000; //
         11'h2ee: return 8'b00000000; //
         11'h2ef: return 8'b00000000; //
         //code x2f
         11'h2f0: return 8'b00000000; //
         11'h2f1: return 8'b00000000; //
         11'h2f2: return 8'b00000000; //
         11'h2f3: return 8'b00000000; //
         11'h2f4: return 8'b00000010; //       *
         11'h2f5: return 8'b00000110; //      **
         11'h2f6: return 8'b00001100; //     **
         11'h2f7: return 8'b00011000; //    **
         11'h2f8: return 8'b00110000; //   **
         11'h2f9: return 8'b01100000; //  **
         11'h2fa: return 8'b11000000; // **
         11'h2fb: return 8'b10000000; // *
         11'h2fc: return 8'b00000000; //
         11'h2fd: return 8'b00000000; //
         11'h2fe: return 8'b00000000; //
         11'h2ff: return 8'b00000000; //
         //code x30
         11'h300: return 8'b00000000; //
         11'h301: return 8'b00000000; //
         11'h302: return 8'b01111100; //  *****
         11'h303: return 8'b11000110; // **   **
         11'h304: return 8'b11000110; // **   **
         11'h305: return 8'b11001110; // **  ***
         11'h306: return 8'b11011110; // ** ****
         11'h307: return 8'b11110110; // **** **
         11'h308: return 8'b11100110; // ***  **
         11'h309: return 8'b11000110; // **   **
         11'h30a: return 8'b11000110; // **   **
         11'h30b: return 8'b01111100; //  *****
         11'h30c: return 8'b00000000; //
         11'h30d: return 8'b00000000; //
         11'h30e: return 8'b00000000; //
         11'h30f: return 8'b00000000; //
         //code x31
         11'h310: return 8'b00000000; //
         11'h311: return 8'b00000000; //
         11'h312: return 8'b00011000; //
         11'h313: return 8'b00111000; //
         11'h314: return 8'b01111000; //    **
         11'h315: return 8'b00011000; //   ***
         11'h316: return 8'b00011000; //  ****
         11'h317: return 8'b00011000; //    **
         11'h318: return 8'b00011000; //    **
         11'h319: return 8'b00011000; //    **
         11'h31a: return 8'b00011000; //    **
         11'h31b: return 8'b01111110; //    **
         11'h31c: return 8'b00000000; //    **
         11'h31d: return 8'b00000000; //  ******
         11'h31e: return 8'b00000000; //
         11'h31f: return 8'b00000000; //
         //code x32
         11'h320: return 8'b00000000; //
         11'h321: return 8'b00000000; //
         11'h322: return 8'b01111100; //  *****
         11'h323: return 8'b11000110; // **   **
         11'h324: return 8'b00000110; //      **
         11'h325: return 8'b00001100; //     **
         11'h326: return 8'b00011000; //    **
         11'h327: return 8'b00110000; //   **
         11'h328: return 8'b01100000; //  **
         11'h329: return 8'b11000000; // **
         11'h32a: return 8'b11000110; // **   **
         11'h32b: return 8'b11111110; // *******
         11'h32c: return 8'b00000000; //
         11'h32d: return 8'b00000000; //
         11'h32e: return 8'b00000000; //
         11'h32f: return 8'b00000000; //
         //code x33
         11'h330: return 8'b00000000; //
         11'h331: return 8'b00000000; //
         11'h332: return 8'b01111100; //  *****
         11'h333: return 8'b11000110; // **   **
         11'h334: return 8'b00000110; //      **
         11'h335: return 8'b00000110; //      **
         11'h336: return 8'b00111100; //   ****
         11'h337: return 8'b00000110; //      **
         11'h338: return 8'b00000110; //      **
         11'h339: return 8'b00000110; //      **
         11'h33a: return 8'b11000110; // **   **
         11'h33b: return 8'b01111100; //  *****
         11'h33c: return 8'b00000000; //
         11'h33d: return 8'b00000000; //
         11'h33e: return 8'b00000000; //
         11'h33f: return 8'b00000000; //
         //code x34
         11'h340: return 8'b00000000; //
         11'h341: return 8'b00000000; //
         11'h342: return 8'b00001100; //     **
         11'h343: return 8'b00011100; //    ***
         11'h344: return 8'b00111100; //   ****
         11'h345: return 8'b01101100; //  ** **
         11'h346: return 8'b11001100; // **  **
         11'h347: return 8'b11111110; // *******
         11'h348: return 8'b00001100; //     **
         11'h349: return 8'b00001100; //     **
         11'h34a: return 8'b00001100; //     **
         11'h34b: return 8'b00011110; //    ****
         11'h34c: return 8'b00000000; //
         11'h34d: return 8'b00000000; //
         11'h34e: return 8'b00000000; //
         11'h34f: return 8'b00000000; //
         //code x35
         11'h350: return 8'b00000000; //
         11'h351: return 8'b00000000; //
         11'h352: return 8'b11111110; // *******
         11'h353: return 8'b11000000; // **
         11'h354: return 8'b11000000; // **
         11'h355: return 8'b11000000; // **
         11'h356: return 8'b11111100; // ******
         11'h357: return 8'b00000110; //      **
         11'h358: return 8'b00000110; //      **
         11'h359: return 8'b00000110; //      **
         11'h35a: return 8'b11000110; // **   **
         11'h35b: return 8'b01111100; //  *****
         11'h35c: return 8'b00000000; //
         11'h35d: return 8'b00000000; //
         11'h35e: return 8'b00000000; //
         11'h35f: return 8'b00000000; //
         //code x36
         11'h360: return 8'b00000000; //
         11'h361: return 8'b00000000; //
         11'h362: return 8'b00111000; //   ***
         11'h363: return 8'b01100000; //  **
         11'h364: return 8'b11000000; // **
         11'h365: return 8'b11000000; // **
         11'h366: return 8'b11111100; // ******
         11'h367: return 8'b11000110; // **   **
         11'h368: return 8'b11000110; // **   **
         11'h369: return 8'b11000110; // **   **
         11'h36a: return 8'b11000110; // **   **
         11'h36b: return 8'b01111100; //  *****
         11'h36c: return 8'b00000000; //
         11'h36d: return 8'b00000000; //
         11'h36e: return 8'b00000000; //
         11'h36f: return 8'b00000000; //
         //code x37
         11'h370: return 8'b00000000; //
         11'h371: return 8'b00000000; //
         11'h372: return 8'b11111110; // *******
         11'h373: return 8'b11000110; // **   **
         11'h374: return 8'b00000110; //      **
         11'h375: return 8'b00000110; //      **
         11'h376: return 8'b00001100; //     **
         11'h377: return 8'b00011000; //    **
         11'h378: return 8'b00110000; //   **
         11'h379: return 8'b00110000; //   **
         11'h37a: return 8'b00110000; //   **
         11'h37b: return 8'b00110000; //   **
         11'h37c: return 8'b00000000; //
         11'h37d: return 8'b00000000; //
         11'h37e: return 8'b00000000; //
         11'h37f: return 8'b00000000; //
         //code x38
         11'h380: return 8'b00000000; //
         11'h381: return 8'b00000000; //
         11'h382: return 8'b01111100; //  *****
         11'h383: return 8'b11000110; // **   **
         11'h384: return 8'b11000110; // **   **
         11'h385: return 8'b11000110; // **   **
         11'h386: return 8'b01111100; //  *****
         11'h387: return 8'b11000110; // **   **
         11'h388: return 8'b11000110; // **   **
         11'h389: return 8'b11000110; // **   **
         11'h38a: return 8'b11000110; // **   **
         11'h38b: return 8'b01111100; //  *****
         11'h38c: return 8'b00000000; //
         11'h38d: return 8'b00000000; //
         11'h38e: return 8'b00000000; //
         11'h38f: return 8'b00000000; //
         //code x39
         11'h390: return 8'b00000000; //
         11'h391: return 8'b00000000; //
         11'h392: return 8'b01111100; //  *****
         11'h393: return 8'b11000110; // **   **
         11'h394: return 8'b11000110; // **   **
         11'h395: return 8'b11000110; // **   **
         11'h396: return 8'b01111110; //  ******
         11'h397: return 8'b00000110; //      **
         11'h398: return 8'b00000110; //      **
         11'h399: return 8'b00000110; //      **
         11'h39a: return 8'b00001100; //     **
         11'h39b: return 8'b01111000; //  ****
         11'h39c: return 8'b00000000; //
         11'h39d: return 8'b00000000; //
         11'h39e: return 8'b00000000; //
         11'h39f: return 8'b00000000; //
         //code x3a
         11'h3a0: return 8'b00000000; //
         11'h3a1: return 8'b00000000; //
         11'h3a2: return 8'b00000000; //
         11'h3a3: return 8'b00000000; //
         11'h3a4: return 8'b00011000; //    **
         11'h3a5: return 8'b00011000; //    **
         11'h3a6: return 8'b00000000; //
         11'h3a7: return 8'b00000000; //
         11'h3a8: return 8'b00000000; //
         11'h3a9: return 8'b00011000; //    **
         11'h3aa: return 8'b00011000; //    **
         11'h3ab: return 8'b00000000; //
         11'h3ac: return 8'b00000000; //
         11'h3ad: return 8'b00000000; //
         11'h3ae: return 8'b00000000; //
         11'h3af: return 8'b00000000; //
         //code x3b
         11'h3b0: return 8'b00000000; //
         11'h3b1: return 8'b00000000; //
         11'h3b2: return 8'b00000000; //
         11'h3b3: return 8'b00000000; //
         11'h3b4: return 8'b00011000; //    **
         11'h3b5: return 8'b00011000; //    **
         11'h3b6: return 8'b00000000; //
         11'h3b7: return 8'b00000000; //
         11'h3b8: return 8'b00000000; //
         11'h3b9: return 8'b00011000; //    **
         11'h3ba: return 8'b00011000; //    **
         11'h3bb: return 8'b00110000; //   **
         11'h3bc: return 8'b00000000; //
         11'h3bd: return 8'b00000000; //
         11'h3be: return 8'b00000000; //
         11'h3bf: return 8'b00000000; //
         //code x3c
         11'h3c0: return 8'b00000000; //
         11'h3c1: return 8'b00000000; //
         11'h3c2: return 8'b00000000; //
         11'h3c3: return 8'b00000110; //      **
         11'h3c4: return 8'b00001100; //     **
         11'h3c5: return 8'b00011000; //    **
         11'h3c6: return 8'b00110000; //   **
         11'h3c7: return 8'b01100000; //  **
         11'h3c8: return 8'b00110000; //   **
         11'h3c9: return 8'b00011000; //    **
         11'h3ca: return 8'b00001100; //     **
         11'h3cb: return 8'b00000110; //      **
         11'h3cc: return 8'b00000000; //
         11'h3cd: return 8'b00000000; //
         11'h3ce: return 8'b00000000; //
         11'h3cf: return 8'b00000000; //
         //code x3d
         11'h3d0: return 8'b00000000; //
         11'h3d1: return 8'b00000000; //
         11'h3d2: return 8'b00000000; //
         11'h3d3: return 8'b00000000; //
         11'h3d4: return 8'b00000000; //
         11'h3d5: return 8'b01111110; //  ******
         11'h3d6: return 8'b00000000; //
         11'h3d7: return 8'b00000000; //
         11'h3d8: return 8'b01111110; //  ******
         11'h3d9: return 8'b00000000; //
         11'h3da: return 8'b00000000; //
         11'h3db: return 8'b00000000; //
         11'h3dc: return 8'b00000000; //
         11'h3dd: return 8'b00000000; //
         11'h3de: return 8'b00000000; //
         11'h3df: return 8'b00000000; //
         //code x3e
         11'h3e0: return 8'b00000000; //
         11'h3e1: return 8'b00000000; //
         11'h3e2: return 8'b00000000; //
         11'h3e3: return 8'b01100000; //  **
         11'h3e4: return 8'b00110000; //   **
         11'h3e5: return 8'b00011000; //    **
         11'h3e6: return 8'b00001100; //     **
         11'h3e7: return 8'b00000110; //      **
         11'h3e8: return 8'b00001100; //     **
         11'h3e9: return 8'b00011000; //    **
         11'h3ea: return 8'b00110000; //   **
         11'h3eb: return 8'b01100000; //  **
         11'h3ec: return 8'b00000000; //
         11'h3ed: return 8'b00000000; //
         11'h3ee: return 8'b00000000; //
         11'h3ef: return 8'b00000000; //
         //code x3f
         11'h3f0: return 8'b00000000; //
         11'h3f1: return 8'b00000000; //
         11'h3f2: return 8'b01111100; //  *****
         11'h3f3: return 8'b11000110; // **   **
         11'h3f4: return 8'b11000110; // **   **
         11'h3f5: return 8'b00001100; //     **
         11'h3f6: return 8'b00011000; //    **
         11'h3f7: return 8'b00011000; //    **
         11'h3f8: return 8'b00011000; //    **
         11'h3f9: return 8'b00000000; //
         11'h3fa: return 8'b00011000; //    **
         11'h3fb: return 8'b00011000; //    **
         11'h3fc: return 8'b00000000; //
         11'h3fd: return 8'b00000000; //
         11'h3fe: return 8'b00000000; //
         11'h3ff: return 8'b00000000; //
        //code x40
         11'h400: return 8'b00000000; //
         11'h401: return 8'b00000000; //
         11'h402: return 8'b01111100; //  *****
         11'h403: return 8'b11000110; // **   **
         11'h404: return 8'b11000110; // **   **
         11'h405: return 8'b11000110; // **   **
         11'h406: return 8'b11011110; // ** ****
         11'h407: return 8'b11011110; // ** ****
         11'h408: return 8'b11011110; // ** ****
         11'h409: return 8'b11011100; // ** ***
         11'h40a: return 8'b11000000; // **
         11'h40b: return 8'b01111100; //  *****
         11'h40c: return 8'b00000000; //
         11'h40d: return 8'b00000000; //
         11'h40e: return 8'b00000000; //
         11'h40f: return 8'b00000000; //
         //code x41
         11'h410: return 8'b00000000; //
         11'h411: return 8'b00000000; //
         11'h412: return 8'b00010000; //    *
         11'h413: return 8'b00111000; //   ***
         11'h414: return 8'b01101100; //  ** **
         11'h415: return 8'b11000110; // **   **
         11'h416: return 8'b11000110; // **   **
         11'h417: return 8'b11111110; // *******
         11'h418: return 8'b11000110; // **   **
         11'h419: return 8'b11000110; // **   **
         11'h41a: return 8'b11000110; // **   **
         11'h41b: return 8'b11000110; // **   **
         11'h41c: return 8'b00000000; //
         11'h41d: return 8'b00000000; //
         11'h41e: return 8'b00000000; //
         11'h41f: return 8'b00000000; //
         //code x42
         11'h420: return 8'b00000000; //
         11'h421: return 8'b00000000; //
         11'h422: return 8'b11111100; // ******
         11'h423: return 8'b01100110; //  **  **
         11'h424: return 8'b01100110; //  **  **
         11'h425: return 8'b01100110; //  **  **
         11'h426: return 8'b01111100; //  *****
         11'h427: return 8'b01100110; //  **  **
         11'h428: return 8'b01100110; //  **  **
         11'h429: return 8'b01100110; //  **  **
         11'h42a: return 8'b01100110; //  **  **
         11'h42b: return 8'b11111100; // ******
         11'h42c: return 8'b00000000; //
         11'h42d: return 8'b00000000; //
         11'h42e: return 8'b00000000; //
         11'h42f: return 8'b00000000; //
         //code x43
         11'h430: return 8'b00000000; //
         11'h431: return 8'b00000000; //
         11'h432: return 8'b00111100; //   ****
         11'h433: return 8'b01100110; //  **  **
         11'h434: return 8'b11000010; // **    *
         11'h435: return 8'b11000000; // **
         11'h436: return 8'b11000000; // **
         11'h437: return 8'b11000000; // **
         11'h438: return 8'b11000000; // **
         11'h439: return 8'b11000010; // **    *
         11'h43a: return 8'b01100110; //  **  **
         11'h43b: return 8'b00111100; //   ****
         11'h43c: return 8'b00000000; //
         11'h43d: return 8'b00000000; //
         11'h43e: return 8'b00000000; //
         11'h43f: return 8'b00000000; //
         //code x44
         11'h440: return 8'b00000000; //
         11'h441: return 8'b00000000; //
         11'h442: return 8'b11111000; // *****
         11'h443: return 8'b01101100; //  ** **
         11'h444: return 8'b01100110; //  **  **
         11'h445: return 8'b01100110; //  **  **
         11'h446: return 8'b01100110; //  **  **
         11'h447: return 8'b01100110; //  **  **
         11'h448: return 8'b01100110; //  **  **
         11'h449: return 8'b01100110; //  **  **
         11'h44a: return 8'b01101100; //  ** **
         11'h44b: return 8'b11111000; // *****
         11'h44c: return 8'b00000000; //
         11'h44d: return 8'b00000000; //
         11'h44e: return 8'b00000000; //
         11'h44f: return 8'b00000000; //
         //code x45
         11'h450: return 8'b00000000; //
         11'h451: return 8'b00000000; //
         11'h452: return 8'b11111110; // *******
         11'h453: return 8'b01100110; //  **  **
         11'h454: return 8'b01100010; //  **   *
         11'h455: return 8'b01101000; //  ** *
         11'h456: return 8'b01111000; //  ****
         11'h457: return 8'b01101000; //  ** *
         11'h458: return 8'b01100000; //  **
         11'h459: return 8'b01100010; //  **   *
         11'h45a: return 8'b01100110; //  **  **
         11'h45b: return 8'b11111110; // *******
         11'h45c: return 8'b00000000; //
         11'h45d: return 8'b00000000; //
         11'h45e: return 8'b00000000; //
         11'h45f: return 8'b00000000; //
         //code x46
         11'h460: return 8'b00000000; //
         11'h461: return 8'b00000000; //
         11'h462: return 8'b11111110; // *******
         11'h463: return 8'b01100110; //  **  **
         11'h464: return 8'b01100010; //  **   *
         11'h465: return 8'b01101000; //  ** *
         11'h466: return 8'b01111000; //  ****
         11'h467: return 8'b01101000; //  ** *
         11'h468: return 8'b01100000; //  **
         11'h469: return 8'b01100000; //  **
         11'h46a: return 8'b01100000; //  **
         11'h46b: return 8'b11110000; // ****
         11'h46c: return 8'b00000000; //
         11'h46d: return 8'b00000000; //
         11'h46e: return 8'b00000000; //
         11'h46f: return 8'b00000000; //
         //code x47
         11'h470: return 8'b00000000; //
         11'h471: return 8'b00000000; //
         11'h472: return 8'b00111100; //   ****
         11'h473: return 8'b01100110; //  **  **
         11'h474: return 8'b11000010; // **    *
         11'h475: return 8'b11000000; // **
         11'h476: return 8'b11000000; // **
         11'h477: return 8'b11011110; // ** ****
         11'h478: return 8'b11000110; // **   **
         11'h479: return 8'b11000110; // **   **
         11'h47a: return 8'b01100110; //  **  **
         11'h47b: return 8'b00111010; //   *** *
         11'h47c: return 8'b00000000; //
         11'h47d: return 8'b00000000; //
         11'h47e: return 8'b00000000; //
         11'h47f: return 8'b00000000; //
         //code x48
         11'h480: return 8'b00000000; //
         11'h481: return 8'b00000000; //
         11'h482: return 8'b11000110; // **   **
         11'h483: return 8'b11000110; // **   **
         11'h484: return 8'b11000110; // **   **
         11'h485: return 8'b11000110; // **   **
         11'h486: return 8'b11111110; // *******
         11'h487: return 8'b11000110; // **   **
         11'h488: return 8'b11000110; // **   **
         11'h489: return 8'b11000110; // **   **
         11'h48a: return 8'b11000110; // **   **
         11'h48b: return 8'b11000110; // **   **
         11'h48c: return 8'b00000000; //
         11'h48d: return 8'b00000000; //
         11'h48e: return 8'b00000000; //
         11'h48f: return 8'b00000000; //
         //code x49
         11'h490: return 8'b00000000; //
         11'h491: return 8'b00000000; //
         11'h492: return 8'b00111100; //   ****
         11'h493: return 8'b00011000; //    **
         11'h494: return 8'b00011000; //    **
         11'h495: return 8'b00011000; //    **
         11'h496: return 8'b00011000; //    **
         11'h497: return 8'b00011000; //    **
         11'h498: return 8'b00011000; //    **
         11'h499: return 8'b00011000; //    **
         11'h49a: return 8'b00011000; //    **
         11'h49b: return 8'b00111100; //   ****
         11'h49c: return 8'b00000000; //
         11'h49d: return 8'b00000000; //
         11'h49e: return 8'b00000000; //
         11'h49f: return 8'b00000000; //
         //code x4a
         11'h4a0: return 8'b00000000; //
         11'h4a1: return 8'b00000000; //
         11'h4a2: return 8'b00011110; //    ****
         11'h4a3: return 8'b00001100; //     **
         11'h4a4: return 8'b00001100; //     **
         11'h4a5: return 8'b00001100; //     **
         11'h4a6: return 8'b00001100; //     **
         11'h4a7: return 8'b00001100; //     **
         11'h4a8: return 8'b11001100; // **  **
         11'h4a9: return 8'b11001100; // **  **
         11'h4aa: return 8'b11001100; // **  **
         11'h4ab: return 8'b01111000; //  ****
         11'h4ac: return 8'b00000000; //
         11'h4ad: return 8'b00000000; //
         11'h4ae: return 8'b00000000; //
         11'h4af: return 8'b00000000; //
         //code x4b
         11'h4b0: return 8'b00000000; //
         11'h4b1: return 8'b00000000; //
         11'h4b2: return 8'b11100110; // ***  **
         11'h4b3: return 8'b01100110; //  **  **
         11'h4b4: return 8'b01100110; //  **  **
         11'h4b5: return 8'b01101100; //  ** **
         11'h4b6: return 8'b01111000; //  ****
         11'h4b7: return 8'b01111000; //  ****
         11'h4b8: return 8'b01101100; //  ** **
         11'h4b9: return 8'b01100110; //  **  **
         11'h4ba: return 8'b01100110; //  **  **
         11'h4bb: return 8'b11100110; // ***  **
         11'h4bc: return 8'b00000000; //
         11'h4bd: return 8'b00000000; //
         11'h4be: return 8'b00000000; //
         11'h4bf: return 8'b00000000; //
         //code x4c
         11'h4c0: return 8'b00000000; //
         11'h4c1: return 8'b00000000; //
         11'h4c2: return 8'b11110000; // ****
         11'h4c3: return 8'b01100000; //  **
         11'h4c4: return 8'b01100000; //  **
         11'h4c5: return 8'b01100000; //  **
         11'h4c6: return 8'b01100000; //  **
         11'h4c7: return 8'b01100000; //  **
         11'h4c8: return 8'b01100000; //  **
         11'h4c9: return 8'b01100010; //  **   *
         11'h4ca: return 8'b01100110; //  **  **
         11'h4cb: return 8'b11111110; // *******
         11'h4cc: return 8'b00000000; //
         11'h4cd: return 8'b00000000; //
         11'h4ce: return 8'b00000000; //
         11'h4cf: return 8'b00000000; //
         //code x4d
         11'h4d0: return 8'b00000000; //
         11'h4d1: return 8'b00000000; //
         11'h4d2: return 8'b11000011; // **    **
         11'h4d3: return 8'b11100111; // ***  ***
         11'h4d4: return 8'b11111111; // ********
         11'h4d5: return 8'b11111111; // ********
         11'h4d6: return 8'b11011011; // ** ** **
         11'h4d7: return 8'b11000011; // **    **
         11'h4d8: return 8'b11000011; // **    **
         11'h4d9: return 8'b11000011; // **    **
         11'h4da: return 8'b11000011; // **    **
         11'h4db: return 8'b11000011; // **    **
         11'h4dc: return 8'b00000000; //
         11'h4dd: return 8'b00000000; //
         11'h4de: return 8'b00000000; //
         11'h4df: return 8'b00000000; //
         //code x4e
         11'h4e0: return 8'b00000000; //
         11'h4e1: return 8'b00000000; //
         11'h4e2: return 8'b11000110; // **   **
         11'h4e3: return 8'b11100110; // ***  **
         11'h4e4: return 8'b11110110; // **** **
         11'h4e5: return 8'b11111110; // *******
         11'h4e6: return 8'b11011110; // ** ****
         11'h4e7: return 8'b11001110; // **  ***
         11'h4e8: return 8'b11000110; // **   **
         11'h4e9: return 8'b11000110; // **   **
         11'h4ea: return 8'b11000110; // **   **
         11'h4eb: return 8'b11000110; // **   **
         11'h4ec: return 8'b00000000; //
         11'h4ed: return 8'b00000000; //
         11'h4ee: return 8'b00000000; //
         11'h4ef: return 8'b00000000; //
         //code x4f
         11'h4f0: return 8'b00000000; //
         11'h4f1: return 8'b00000000; //
         11'h4f2: return 8'b01111100; //  *****
         11'h4f3: return 8'b11000110; // **   **
         11'h4f4: return 8'b11000110; // **   **
         11'h4f5: return 8'b11000110; // **   **
         11'h4f6: return 8'b11000110; // **   **
         11'h4f7: return 8'b11000110; // **   **
         11'h4f8: return 8'b11000110; // **   **
         11'h4f9: return 8'b11000110; // **   **
         11'h4fa: return 8'b11000110; // **   **
         11'h4fb: return 8'b01111100; //  *****
         11'h4fc: return 8'b00000000; //
         11'h4fd: return 8'b00000000; //
         11'h4fe: return 8'b00000000; //
         11'h4ff: return 8'b00000000; //
         //code x50
         11'h500: return 8'b00000000; //
         11'h501: return 8'b00000000; //
         11'h502: return 8'b11111100; // ******
         11'h503: return 8'b01100110; //  **  **
         11'h504: return 8'b01100110; //  **  **
         11'h505: return 8'b01100110; //  **  **
         11'h506: return 8'b01111100; //  *****
         11'h507: return 8'b01100000; //  **
         11'h508: return 8'b01100000; //  **
         11'h509: return 8'b01100000; //  **
         11'h50a: return 8'b01100000; //  **
         11'h50b: return 8'b11110000; // ****
         11'h50c: return 8'b00000000; //
         11'h50d: return 8'b00000000; //
         11'h50e: return 8'b00000000; //
         11'h50f: return 8'b00000000; //
         //code x510f
         11'h510: return 8'b00000000; //
         11'h511: return 8'b00000000; //
         11'h512: return 8'b01111100; //  *****
         11'h513: return 8'b11000110; // **   **
         11'h514: return 8'b11000110; // **   **
         11'h515: return 8'b11000110; // **   **
         11'h516: return 8'b11000110; // **   **
         11'h517: return 8'b11000110; // **   **
         11'h518: return 8'b11000110; // **   **
         11'h519: return 8'b11010110; // ** * **
         11'h51a: return 8'b11011110; // ** ****
         11'h51b: return 8'b01111100; //  *****
         11'h51c: return 8'b00001100; //     **
         11'h51d: return 8'b00001110; //     ***
         11'h51e: return 8'b00000000; //
         11'h51f: return 8'b00000000; //
         //code x52
         11'h520: return 8'b00000000; //
         11'h521: return 8'b00000000; //
         11'h522: return 8'b11111100; // ******
         11'h523: return 8'b01100110; //  **  **
         11'h524: return 8'b01100110; //  **  **
         11'h525: return 8'b01100110; //  **  **
         11'h526: return 8'b01111100; //  *****
         11'h527: return 8'b01101100; //  ** **
         11'h528: return 8'b01100110; //  **  **
         11'h529: return 8'b01100110; //  **  **
         11'h52a: return 8'b01100110; //  **  **
         11'h52b: return 8'b11100110; // ***  **
         11'h52c: return 8'b00000000; //
         11'h52d: return 8'b00000000; //
         11'h52e: return 8'b00000000; //
         11'h52f: return 8'b00000000; //
         //code x53
         11'h530: return 8'b00000000; //
         11'h531: return 8'b00000000; //
         11'h532: return 8'b01111100; //  *****
         11'h533: return 8'b11000110; // **   **
         11'h534: return 8'b11000110; // **   **
         11'h535: return 8'b01100000; //  **
         11'h536: return 8'b00111000; //   ***
         11'h537: return 8'b00001100; //     **
         11'h538: return 8'b00000110; //      **
         11'h539: return 8'b11000110; // **   **
         11'h53a: return 8'b11000110; // **   **
         11'h53b: return 8'b01111100; //  *****
         11'h53c: return 8'b00000000; //
         11'h53d: return 8'b00000000; //
         11'h53e: return 8'b00000000; //
         11'h53f: return 8'b00000000; //
         //code x54
         11'h540: return 8'b00000000; //
         11'h541: return 8'b00000000; //
         11'h542: return 8'b11111111; // ********
         11'h543: return 8'b11011011; // ** ** **
         11'h544: return 8'b10011001; // *  **  *
         11'h545: return 8'b00011000; //    **
         11'h546: return 8'b00011000; //    **
         11'h547: return 8'b00011000; //    **
         11'h548: return 8'b00011000; //    **
         11'h549: return 8'b00011000; //    **
         11'h54a: return 8'b00011000; //    **
         11'h54b: return 8'b00111100; //   ****
         11'h54c: return 8'b00000000; //
         11'h54d: return 8'b00000000; //
         11'h54e: return 8'b00000000; //
         11'h54f: return 8'b00000000; //
         //code x55
         11'h550: return 8'b00000000; //
         11'h551: return 8'b00000000; //
         11'h552: return 8'b11000110; // **   **
         11'h553: return 8'b11000110; // **   **
         11'h554: return 8'b11000110; // **   **
         11'h555: return 8'b11000110; // **   **
         11'h556: return 8'b11000110; // **   **
         11'h557: return 8'b11000110; // **   **
         11'h558: return 8'b11000110; // **   **
         11'h559: return 8'b11000110; // **   **
         11'h55a: return 8'b11000110; // **   **
         11'h55b: return 8'b01111100; //  *****
         11'h55c: return 8'b00000000; //
         11'h55d: return 8'b00000000; //
         11'h55e: return 8'b00000000; //
         11'h55f: return 8'b00000000; //
         //code x56
         11'h560: return 8'b00000000; //
         11'h561: return 8'b00000000; //
         11'h562: return 8'b11000011; // **    **
         11'h563: return 8'b11000011; // **    **
         11'h564: return 8'b11000011; // **    **
         11'h565: return 8'b11000011; // **    **
         11'h566: return 8'b11000011; // **    **
         11'h567: return 8'b11000011; // **    **
         11'h568: return 8'b11000011; // **    **
         11'h569: return 8'b01100110; //  **  **
         11'h56a: return 8'b00111100; //   ****
         11'h56b: return 8'b00011000; //    **
         11'h56c: return 8'b00000000; //
         11'h56d: return 8'b00000000; //
         11'h56e: return 8'b00000000; //
         11'h56f: return 8'b00000000; //
         //code x57
         11'h570: return 8'b00000000; //
         11'h571: return 8'b00000000; //
         11'h572: return 8'b11000011; // **    **
         11'h573: return 8'b11000011; // **    **
         11'h574: return 8'b11000011; // **    **
         11'h575: return 8'b11000011; // **    **
         11'h576: return 8'b11000011; // **    **
         11'h577: return 8'b11011011; // ** ** **
         11'h578: return 8'b11011011; // ** ** **
         11'h579: return 8'b11111111; // ********
         11'h57a: return 8'b01100110; //  **  **
         11'h57b: return 8'b01100110; //  **  **
         11'h57c: return 8'b00000000; //
         11'h57d: return 8'b00000000; //
         11'h57e: return 8'b00000000; //
         11'h57f: return 8'b00000000; //
         //code x58
         11'h580: return 8'b00000000; //
         11'h581: return 8'b00000000; //
         11'h582: return 8'b11000011; // **    **
         11'h583: return 8'b11000011; // **    **
         11'h584: return 8'b01100110; //  **  **
         11'h585: return 8'b00111100; //   ****
         11'h586: return 8'b00011000; //    **
         11'h587: return 8'b00011000; //    **
         11'h588: return 8'b00111100; //   ****
         11'h589: return 8'b01100110; //  **  **
         11'h58a: return 8'b11000011; // **    **
         11'h58b: return 8'b11000011; // **    **
         11'h58c: return 8'b00000000; //
         11'h58d: return 8'b00000000; //
         11'h58e: return 8'b00000000; //
         11'h58f: return 8'b00000000; //
         //code x59
         11'h590: return 8'b00000000; //
         11'h591: return 8'b00000000; //
         11'h592: return 8'b11000011; // **    **
         11'h593: return 8'b11000011; // **    **
         11'h594: return 8'b11000011; // **    **
         11'h595: return 8'b01100110; //  **  **
         11'h596: return 8'b00111100; //   ****
         11'h597: return 8'b00011000; //    **
         11'h598: return 8'b00011000; //    **
         11'h599: return 8'b00011000; //    **
         11'h59a: return 8'b00011000; //    **
         11'h59b: return 8'b00111100; //   ****
         11'h59c: return 8'b00000000; //
         11'h59d: return 8'b00000000; //
         11'h59e: return 8'b00000000; //
         11'h59f: return 8'b00000000; //
         //code x5a
         11'h5a0: return 8'b00000000; //
         11'h5a1: return 8'b00000000; //
         11'h5a2: return 8'b11111111; // ********
         11'h5a3: return 8'b11000011; // **    **
         11'h5a4: return 8'b10000110; // *    **
         11'h5a5: return 8'b00001100; //     **
         11'h5a6: return 8'b00011000; //    **
         11'h5a7: return 8'b00110000; //   **
         11'h5a8: return 8'b01100000; //  **
         11'h5a9: return 8'b11000001; // **     *
         11'h5aa: return 8'b11000011; // **    **
         11'h5ab: return 8'b11111111; // ********
         11'h5ac: return 8'b00000000; //
         11'h5ad: return 8'b00000000; //
         11'h5ae: return 8'b00000000; //
         11'h5af: return 8'b00000000; //
         //code x5b
         11'h5b0: return 8'b00000000; //
         11'h5b1: return 8'b00000000; //
         11'h5b2: return 8'b00111100; //   ****
         11'h5b3: return 8'b00110000; //   **
         11'h5b4: return 8'b00110000; //   **
         11'h5b5: return 8'b00110000; //   **
         11'h5b6: return 8'b00110000; //   **
         11'h5b7: return 8'b00110000; //   **
         11'h5b8: return 8'b00110000; //   **
         11'h5b9: return 8'b00110000; //   **
         11'h5ba: return 8'b00110000; //   **
         11'h5bb: return 8'b00111100; //   ****
         11'h5bc: return 8'b00000000; //
         11'h5bd: return 8'b00000000; //
         11'h5be: return 8'b00000000; //
         11'h5bf: return 8'b00000000; //
         //code x5c
         11'h5c0: return 8'b00000000; //
         11'h5c1: return 8'b00000000; //
         11'h5c2: return 8'b00000000; //
         11'h5c3: return 8'b10000000; // *
         11'h5c4: return 8'b11000000; // **
         11'h5c5: return 8'b11100000; // ***
         11'h5c6: return 8'b01110000; //  ***
         11'h5c7: return 8'b00111000; //   ***
         11'h5c8: return 8'b00011100; //    ***
         11'h5c9: return 8'b00001110; //     ***
         11'h5ca: return 8'b00000110; //      **
         11'h5cb: return 8'b00000010; //       *
         11'h5cc: return 8'b00000000; //
         11'h5cd: return 8'b00000000; //
         11'h5ce: return 8'b00000000; //
         11'h5cf: return 8'b00000000; //
         //code x5d
         11'h5d0: return 8'b00000000; //
         11'h5d1: return 8'b00000000; //
         11'h5d2: return 8'b00111100; //   ****
         11'h5d3: return 8'b00001100; //     **
         11'h5d4: return 8'b00001100; //     **
         11'h5d5: return 8'b00001100; //     **
         11'h5d6: return 8'b00001100; //     **
         11'h5d7: return 8'b00001100; //     **
         11'h5d8: return 8'b00001100; //     **
         11'h5d9: return 8'b00001100; //     **
         11'h5da: return 8'b00001100; //     **
         11'h5db: return 8'b00111100; //   ****
         11'h5dc: return 8'b00000000; //
         11'h5dd: return 8'b00000000; //
         11'h5de: return 8'b00000000; //
         11'h5df: return 8'b00000000; //
         //code x5e
         11'h5e0: return 8'b00010000; //    *
         11'h5e1: return 8'b00111000; //   ***
         11'h5e2: return 8'b01101100; //  ** **
         11'h5e3: return 8'b11000110; // **   **
         11'h5e4: return 8'b00000000; //
         11'h5e5: return 8'b00000000; //
         11'h5e6: return 8'b00000000; //
         11'h5e7: return 8'b00000000; //
         11'h5e8: return 8'b00000000; //
         11'h5e9: return 8'b00000000; //
         11'h5ea: return 8'b00000000; //
         11'h5eb: return 8'b00000000; //
         11'h5ec: return 8'b00000000; //
         11'h5ed: return 8'b00000000; //
         11'h5ee: return 8'b00000000; //
         11'h5ef: return 8'b00000000; //
         //code x5f
         11'h5f0: return 8'b00000000; //
         11'h5f1: return 8'b00000000; //
         11'h5f2: return 8'b00000000; //
         11'h5f3: return 8'b00000000; //
         11'h5f4: return 8'b00000000; //
         11'h5f5: return 8'b00000000; //
         11'h5f6: return 8'b00000000; //
         11'h5f7: return 8'b00000000; //
         11'h5f8: return 8'b00000000; //
         11'h5f9: return 8'b00000000; //
         11'h5fa: return 8'b00000000; //
         11'h5fb: return 8'b00000000; //
         11'h5fc: return 8'b00000000; //
         11'h5fd: return 8'b11111111; // ********
         11'h5fe: return 8'b00000000; //
         11'h5ff: return 8'b00000000; //
         //code x60
         11'h600: return 8'b00110000; //   **
         11'h601: return 8'b00110000; //   **
         11'h602: return 8'b00011000; //    **
         11'h603: return 8'b00000000; //
         11'h604: return 8'b00000000; //
         11'h605: return 8'b00000000; //
         11'h606: return 8'b00000000; //
         11'h607: return 8'b00000000; //
         11'h608: return 8'b00000000; //
         11'h609: return 8'b00000000; //
         11'h60a: return 8'b00000000; //
         11'h60b: return 8'b00000000; //
         11'h60c: return 8'b00000000; //
         11'h60d: return 8'b00000000; //
         11'h60e: return 8'b00000000; //
         11'h60f: return 8'b00000000; //
         //code x61
         11'h610: return 8'b00000000; //
         11'h611: return 8'b00000000; //
         11'h612: return 8'b00000000; //
         11'h613: return 8'b00000000; //
         11'h614: return 8'b00000000; //
         11'h615: return 8'b01111000; //  ****
         11'h616: return 8'b00001100; //     **
         11'h617: return 8'b01111100; //  *****
         11'h618: return 8'b11001100; // **  **
         11'h619: return 8'b11001100; // **  **
         11'h61a: return 8'b11001100; // **  **
         11'h61b: return 8'b01110110; //  *** **
         11'h61c: return 8'b00000000; //
         11'h61d: return 8'b00000000; //
         11'h61e: return 8'b00000000; //
         11'h61f: return 8'b00000000; //
         //code x62
         11'h620: return 8'b00000000; //
         11'h621: return 8'b00000000; //
         11'h622: return 8'b11100000; //  ***
         11'h623: return 8'b01100000; //   **
         11'h624: return 8'b01100000; //   **
         11'h625: return 8'b01111000; //   ****
         11'h626: return 8'b01101100; //   ** **
         11'h627: return 8'b01100110; //   **  **
         11'h628: return 8'b01100110; //   **  **
         11'h629: return 8'b01100110; //   **  **
         11'h62a: return 8'b01100110; //   **  **
         11'h62b: return 8'b01111100; //   *****
         11'h62c: return 8'b00000000; //
         11'h62d: return 8'b00000000; //
         11'h62e: return 8'b00000000; //
         11'h62f: return 8'b00000000; //
         //code x63
         11'h630: return 8'b00000000; //
         11'h631: return 8'b00000000; //
         11'h632: return 8'b00000000; //
         11'h633: return 8'b00000000; //
         11'h634: return 8'b00000000; //
         11'h635: return 8'b01111100; //  *****
         11'h636: return 8'b11000110; // **   **
         11'h637: return 8'b11000000; // **
         11'h638: return 8'b11000000; // **
         11'h639: return 8'b11000000; // **
         11'h63a: return 8'b11000110; // **   **
         11'h63b: return 8'b01111100; //  *****
         11'h63c: return 8'b00000000; //
         11'h63d: return 8'b00000000; //
         11'h63e: return 8'b00000000; //
         11'h63f: return 8'b00000000; //
         //code x64
         11'h640: return 8'b00000000; //
         11'h641: return 8'b00000000; //
         11'h642: return 8'b00011100; //    ***
         11'h643: return 8'b00001100; //     **
         11'h644: return 8'b00001100; //     **
         11'h645: return 8'b00111100; //   ****
         11'h646: return 8'b01101100; //  ** **
         11'h647: return 8'b11001100; // **  **
         11'h648: return 8'b11001100; // **  **
         11'h649: return 8'b11001100; // **  **
         11'h64a: return 8'b11001100; // **  **
         11'h64b: return 8'b01110110; //  *** **
         11'h64c: return 8'b00000000; //
         11'h64d: return 8'b00000000; //
         11'h64e: return 8'b00000000; //
         11'h64f: return 8'b00000000; //
         //code x65
         11'h650: return 8'b00000000; //
         11'h651: return 8'b00000000; //
         11'h652: return 8'b00000000; //
         11'h653: return 8'b00000000; //
         11'h654: return 8'b00000000; //
         11'h655: return 8'b01111100; //  *****
         11'h656: return 8'b11000110; // **   **
         11'h657: return 8'b11111110; // *******
         11'h658: return 8'b11000000; // **
         11'h659: return 8'b11000000; // **
         11'h65a: return 8'b11000110; // **   **
         11'h65b: return 8'b01111100; //  *****
         11'h65c: return 8'b00000000; //
         11'h65d: return 8'b00000000; //
         11'h65e: return 8'b00000000; //
         11'h65f: return 8'b00000000; //
         //code x66
         11'h660: return 8'b00000000; //
         11'h661: return 8'b00000000; //
         11'h662: return 8'b00111000; //   ***
         11'h663: return 8'b01101100; //  ** **
         11'h664: return 8'b01100100; //  **  *
         11'h665: return 8'b01100000; //  **
         11'h666: return 8'b11110000; // ****
         11'h667: return 8'b01100000; //  **
         11'h668: return 8'b01100000; //  **
         11'h669: return 8'b01100000; //  **
         11'h66a: return 8'b01100000; //  **
         11'h66b: return 8'b11110000; // ****
         11'h66c: return 8'b00000000; //
         11'h66d: return 8'b00000000; //
         11'h66e: return 8'b00000000; //
         11'h66f: return 8'b00000000; //
         //code x67
         11'h670: return 8'b00000000; //
         11'h671: return 8'b00000000; //
         11'h672: return 8'b00000000; //
         11'h673: return 8'b00000000; //
         11'h674: return 8'b00000000; //
         11'h675: return 8'b01110110; //  *** **
         11'h676: return 8'b11001100; // **  **
         11'h677: return 8'b11001100; // **  **
         11'h678: return 8'b11001100; // **  **
         11'h679: return 8'b11001100; // **  **
         11'h67a: return 8'b11001100; // **  **
         11'h67b: return 8'b01111100; //  *****
         11'h67c: return 8'b00001100; //     **
         11'h67d: return 8'b11001100; // **  **
         11'h67e: return 8'b01111000; //  ****
         11'h67f: return 8'b00000000; //
         //code x68
         11'h680: return 8'b00000000; //
         11'h681: return 8'b00000000; //
         11'h682: return 8'b11100000; // ***
         11'h683: return 8'b01100000; //  **
         11'h684: return 8'b01100000; //  **
         11'h685: return 8'b01101100; //  ** **
         11'h686: return 8'b01110110; //  *** **
         11'h687: return 8'b01100110; //  **  **
         11'h688: return 8'b01100110; //  **  **
         11'h689: return 8'b01100110; //  **  **
         11'h68a: return 8'b01100110; //  **  **
         11'h68b: return 8'b11100110; // ***  **
         11'h68c: return 8'b00000000; //
         11'h68d: return 8'b00000000; //
         11'h68e: return 8'b00000000; //
         11'h68f: return 8'b00000000; //
         //code x69
         11'h690: return 8'b00000000; //
         11'h691: return 8'b00000000; //
         11'h692: return 8'b00011000; //    **
         11'h693: return 8'b00011000; //    **
         11'h694: return 8'b00000000; //
         11'h695: return 8'b00111000; //   ***
         11'h696: return 8'b00011000; //    **
         11'h697: return 8'b00011000; //    **
         11'h698: return 8'b00011000; //    **
         11'h699: return 8'b00011000; //    **
         11'h69a: return 8'b00011000; //    **
         11'h69b: return 8'b00111100; //   ****
         11'h69c: return 8'b00000000; //
         11'h69d: return 8'b00000000; //
         11'h69e: return 8'b00000000; //
         11'h69f: return 8'b00000000; //
         //code x6a
         11'h6a0: return 8'b00000000; //
         11'h6a1: return 8'b00000000; //
         11'h6a2: return 8'b00000110; //      **
         11'h6a3: return 8'b00000110; //      **
         11'h6a4: return 8'b00000000; //
         11'h6a5: return 8'b00001110; //     ***
         11'h6a6: return 8'b00000110; //      **
         11'h6a7: return 8'b00000110; //      **
         11'h6a8: return 8'b00000110; //      **
         11'h6a9: return 8'b00000110; //      **
         11'h6aa: return 8'b00000110; //      **
         11'h6ab: return 8'b00000110; //      **
         11'h6ac: return 8'b01100110; //  **  **
         11'h6ad: return 8'b01100110; //  **  **
         11'h6ae: return 8'b00111100; //   ****
         11'h6af: return 8'b00000000; //
         //code x6b
         11'h6b0: return 8'b00000000; //
         11'h6b1: return 8'b00000000; //
         11'h6b2: return 8'b11100000; // ***
         11'h6b3: return 8'b01100000; //  **
         11'h6b4: return 8'b01100000; //  **
         11'h6b5: return 8'b01100110; //  **  **
         11'h6b6: return 8'b01101100; //  ** **
         11'h6b7: return 8'b01111000; //  ****
         11'h6b8: return 8'b01111000; //  ****
         11'h6b9: return 8'b01101100; //  ** **
         11'h6ba: return 8'b01100110; //  **  **
         11'h6bb: return 8'b11100110; // ***  **
         11'h6bc: return 8'b00000000; //
         11'h6bd: return 8'b00000000; //
         11'h6be: return 8'b00000000; //
         11'h6bf: return 8'b00000000; //
         //code x6c
         11'h6c0: return 8'b00000000; //
         11'h6c1: return 8'b00000000; //
         11'h6c2: return 8'b00111000; //   ***
         11'h6c3: return 8'b00011000; //    **
         11'h6c4: return 8'b00011000; //    **
         11'h6c5: return 8'b00011000; //    **
         11'h6c6: return 8'b00011000; //    **
         11'h6c7: return 8'b00011000; //    **
         11'h6c8: return 8'b00011000; //    **
         11'h6c9: return 8'b00011000; //    **
         11'h6ca: return 8'b00011000; //    **
         11'h6cb: return 8'b00111100; //   ****
         11'h6cc: return 8'b00000000; //
         11'h6cd: return 8'b00000000; //
         11'h6ce: return 8'b00000000; //
         11'h6cf: return 8'b00000000; //
         //code x6d
         11'h6d0: return 8'b00000000; //
         11'h6d1: return 8'b00000000; //
         11'h6d2: return 8'b00000000; //
         11'h6d3: return 8'b00000000; //
         11'h6d4: return 8'b00000000; //
         11'h6d5: return 8'b11100110; // ***  **
         11'h6d6: return 8'b11111111; // ********
         11'h6d7: return 8'b11011011; // ** ** **
         11'h6d8: return 8'b11011011; // ** ** **
         11'h6d9: return 8'b11011011; // ** ** **
         11'h6da: return 8'b11011011; // ** ** **
         11'h6db: return 8'b11011011; // ** ** **
         11'h6dc: return 8'b00000000; //
         11'h6dd: return 8'b00000000; //
         11'h6de: return 8'b00000000; //
         11'h6df: return 8'b00000000; //
         //code x6e
         11'h6e0: return 8'b00000000; //
         11'h6e1: return 8'b00000000; //
         11'h6e2: return 8'b00000000; //
         11'h6e3: return 8'b00000000; //
         11'h6e4: return 8'b00000000; //
         11'h6e5: return 8'b11011100; // ** ***
         11'h6e6: return 8'b01100110; //  **  **
         11'h6e7: return 8'b01100110; //  **  **
         11'h6e8: return 8'b01100110; //  **  **
         11'h6e9: return 8'b01100110; //  **  **
         11'h6ea: return 8'b01100110; //  **  **
         11'h6eb: return 8'b01100110; //  **  **
         11'h6ec: return 8'b00000000; //
         11'h6ed: return 8'b00000000; //
         11'h6ee: return 8'b00000000; //
         11'h6ef: return 8'b00000000; //
         //code x6f
         11'h6f0: return 8'b00000000; //
         11'h6f1: return 8'b00000000; //
         11'h6f2: return 8'b00000000; //
         11'h6f3: return 8'b00000000; //
         11'h6f4: return 8'b00000000; //
         11'h6f5: return 8'b01111100; //  *****
         11'h6f6: return 8'b11000110; // **   **
         11'h6f7: return 8'b11000110; // **   **
         11'h6f8: return 8'b11000110; // **   **
         11'h6f9: return 8'b11000110; // **   **
         11'h6fa: return 8'b11000110; // **   **
         11'h6fb: return 8'b01111100; //  *****
         11'h6fc: return 8'b00000000; //
         11'h6fd: return 8'b00000000; //
         11'h6fe: return 8'b00000000; //
         11'h6ff: return 8'b00000000; //
         //code x70
         11'h700: return 8'b00000000; //
         11'h701: return 8'b00000000; //
         11'h702: return 8'b00000000; //
         11'h703: return 8'b00000000; //
         11'h704: return 8'b00000000; //
         11'h705: return 8'b11011100; // ** ***
         11'h706: return 8'b01100110; //  **  **
         11'h707: return 8'b01100110; //  **  **
         11'h708: return 8'b01100110; //  **  **
         11'h709: return 8'b01100110; //  **  **
         11'h70a: return 8'b01100110; //  **  **
         11'h70b: return 8'b01111100; //  *****
         11'h70c: return 8'b01100000; //  **
         11'h70d: return 8'b01100000; //  **
         11'h70e: return 8'b11110000; // ****
         11'h70f: return 8'b00000000; //
         //code x71
         11'h710: return 8'b00000000; //
         11'h711: return 8'b00000000; //
         11'h712: return 8'b00000000; //
         11'h713: return 8'b00000000; //
         11'h714: return 8'b00000000; //
         11'h715: return 8'b01110110; //  *** **
         11'h716: return 8'b11001100; // **  **
         11'h717: return 8'b11001100; // **  **
         11'h718: return 8'b11001100; // **  **
         11'h719: return 8'b11001100; // **  **
         11'h71a: return 8'b11001100; // **  **
         11'h71b: return 8'b01111100; //  *****
         11'h71c: return 8'b00001100; //     **
         11'h71d: return 8'b00001100; //     **
         11'h71e: return 8'b00011110; //    ****
         11'h71f: return 8'b00000000; //
         //code x72
         11'h720: return 8'b00000000; //
         11'h721: return 8'b00000000; //
         11'h722: return 8'b00000000; //
         11'h723: return 8'b00000000; //
         11'h724: return 8'b00000000; //
         11'h725: return 8'b11011100; // ** ***
         11'h726: return 8'b01110110; //  *** **
         11'h727: return 8'b01100110; //  **  **
         11'h728: return 8'b01100000; //  **
         11'h729: return 8'b01100000; //  **
         11'h72a: return 8'b01100000; //  **
         11'h72b: return 8'b11110000; // ****
         11'h72c: return 8'b00000000; //
         11'h72d: return 8'b00000000; //
         11'h72e: return 8'b00000000; //
         11'h72f: return 8'b00000000; //
         //code x73
         11'h730: return 8'b00000000; //
         11'h731: return 8'b00000000; //
         11'h732: return 8'b00000000; //
         11'h733: return 8'b00000000; //
         11'h734: return 8'b00000000; //
         11'h735: return 8'b01111100; //  *****
         11'h736: return 8'b11000110; // **   **
         11'h737: return 8'b01100000; //  **
         11'h738: return 8'b00111000; //   ***
         11'h739: return 8'b00001100; //     **
         11'h73a: return 8'b11000110; // **   **
         11'h73b: return 8'b01111100; //  *****
         11'h73c: return 8'b00000000; //
         11'h73d: return 8'b00000000; //
         11'h73e: return 8'b00000000; //
         11'h73f: return 8'b00000000; //
         //code x74
         11'h740: return 8'b00000000; //
         11'h741: return 8'b00000000; //
         11'h742: return 8'b00010000; //    *
         11'h743: return 8'b00110000; //   **
         11'h744: return 8'b00110000; //   **
         11'h745: return 8'b11111100; // ******
         11'h746: return 8'b00110000; //   **
         11'h747: return 8'b00110000; //   **
         11'h748: return 8'b00110000; //   **
         11'h749: return 8'b00110000; //   **
         11'h74a: return 8'b00110110; //   ** **
         11'h74b: return 8'b00011100; //    ***
         11'h74c: return 8'b00000000; //
         11'h74d: return 8'b00000000; //
         11'h74e: return 8'b00000000; //
         11'h74f: return 8'b00000000; //
         //code x75
         11'h750: return 8'b00000000; //
         11'h751: return 8'b00000000; //
         11'h752: return 8'b00000000; //
         11'h753: return 8'b00000000; //
         11'h754: return 8'b00000000; //
         11'h755: return 8'b11001100; // **  **
         11'h756: return 8'b11001100; // **  **
         11'h757: return 8'b11001100; // **  **
         11'h758: return 8'b11001100; // **  **
         11'h759: return 8'b11001100; // **  **
         11'h75a: return 8'b11001100; // **  **
         11'h75b: return 8'b01110110; //  *** **
         11'h75c: return 8'b00000000; //
         11'h75d: return 8'b00000000; //
         11'h75e: return 8'b00000000; //
         11'h75f: return 8'b00000000; //
         //code x76
         11'h760: return 8'b00000000; //
         11'h761: return 8'b00000000; //
         11'h762: return 8'b00000000; //
         11'h763: return 8'b00000000; //
         11'h764: return 8'b00000000; //
         11'h765: return 8'b11000011; // **    **
         11'h766: return 8'b11000011; // **    **
         11'h767: return 8'b11000011; // **    **
         11'h768: return 8'b11000011; // **    **
         11'h769: return 8'b01100110; //  **  **
         11'h76a: return 8'b00111100; //   ****
         11'h76b: return 8'b00011000; //    **
         11'h76c: return 8'b00000000; //
         11'h76d: return 8'b00000000; //
         11'h76e: return 8'b00000000; //
         11'h76f: return 8'b00000000; //
         //code x77
         11'h770: return 8'b00000000; //
         11'h771: return 8'b00000000; //
         11'h772: return 8'b00000000; //
         11'h773: return 8'b00000000; //
         11'h774: return 8'b00000000; //
         11'h775: return 8'b11000011; // **    **
         11'h776: return 8'b11000011; // **    **
         11'h777: return 8'b11000011; // **    **
         11'h778: return 8'b11011011; // ** ** **
         11'h779: return 8'b11011011; // ** ** **
         11'h77a: return 8'b11111111; // ********
         11'h77b: return 8'b01100110; //  **  **
         11'h77c: return 8'b00000000; //
         11'h77d: return 8'b00000000; //
         11'h77e: return 8'b00000000; //
         11'h77f: return 8'b00000000; //
         //code x78
         11'h780: return 8'b00000000; //
         11'h781: return 8'b00000000; //
         11'h782: return 8'b00000000; //
         11'h783: return 8'b00000000; //
         11'h784: return 8'b00000000; //
         11'h785: return 8'b11000011; // **    **
         11'h786: return 8'b01100110; //  **  **
         11'h787: return 8'b00111100; //   ****
         11'h788: return 8'b00011000; //    **
         11'h789: return 8'b00111100; //   ****
         11'h78a: return 8'b01100110; //  **  **
         11'h78b: return 8'b11000011; // **    **
         11'h78c: return 8'b00000000; //
         11'h78d: return 8'b00000000; //
         11'h78e: return 8'b00000000; //
         11'h78f: return 8'b00000000; //
         //code x79
         11'h790: return 8'b00000000; //
         11'h791: return 8'b00000000; //
         11'h792: return 8'b00000000; //
         11'h793: return 8'b00000000; //
         11'h794: return 8'b00000000; //
         11'h795: return 8'b11000110; // **   **
         11'h796: return 8'b11000110; // **   **
         11'h797: return 8'b11000110; // **   **
         11'h798: return 8'b11000110; // **   **
         11'h799: return 8'b11000110; // **   **
         11'h79a: return 8'b11000110; // **   **
         11'h79b: return 8'b01111110; //  ******
         11'h79c: return 8'b00000110; //      **
         11'h79d: return 8'b00001100; //     **
         11'h79e: return 8'b11111000; // *****
         11'h79f: return 8'b00000000; //
         //code x7a
         11'h7a0: return 8'b00000000; //
         11'h7a1: return 8'b00000000; //
         11'h7a2: return 8'b00000000; //
         11'h7a3: return 8'b00000000; //
         11'h7a4: return 8'b00000000; //
         11'h7a5: return 8'b11111110; // *******
         11'h7a6: return 8'b11001100; // **  **
         11'h7a7: return 8'b00011000; //    **
         11'h7a8: return 8'b00110000; //   **
         11'h7a9: return 8'b01100000; //  **
         11'h7aa: return 8'b11000110; // **   **
         11'h7ab: return 8'b11111110; // *******
         11'h7ac: return 8'b00000000; //
         11'h7ad: return 8'b00000000; //
         11'h7ae: return 8'b00000000; //
         11'h7af: return 8'b00000000; //
         //code x7b
         11'h7b0: return 8'b00000000; //
         11'h7b1: return 8'b00000000; //
         11'h7b2: return 8'b00001110; //     ***
         11'h7b3: return 8'b00011000; //    **
         11'h7b4: return 8'b00011000; //    **
         11'h7b5: return 8'b00011000; //    **
         11'h7b6: return 8'b01110000; //  ***
         11'h7b7: return 8'b00011000; //    **
         11'h7b8: return 8'b00011000; //    **
         11'h7b9: return 8'b00011000; //    **
         11'h7ba: return 8'b00011000; //    **
         11'h7bb: return 8'b00001110; //     ***
         11'h7bc: return 8'b00000000; //
         11'h7bd: return 8'b00000000; //
         11'h7be: return 8'b00000000; //
         11'h7bf: return 8'b00000000; //
         //code x7c
         11'h7c0: return 8'b00000000; //
         11'h7c1: return 8'b00000000; //
         11'h7c2: return 8'b00011000; //    **
         11'h7c3: return 8'b00011000; //    **
         11'h7c4: return 8'b00011000; //    **
         11'h7c5: return 8'b00011000; //    **
         11'h7c6: return 8'b00000000; //
         11'h7c7: return 8'b00011000; //    **
         11'h7c8: return 8'b00011000; //    **
         11'h7c9: return 8'b00011000; //    **
         11'h7ca: return 8'b00011000; //    **
         11'h7cb: return 8'b00011000; //    **
         11'h7cc: return 8'b00000000; //
         11'h7cd: return 8'b00000000; //
         11'h7ce: return 8'b00000000; //
         11'h7cf: return 8'b00000000; //
         //code x7d
         11'h7d0: return 8'b00000000; //
         11'h7d1: return 8'b00000000; //
         11'h7d2: return 8'b01110000; //  ***
         11'h7d3: return 8'b00011000; //    **
         11'h7d4: return 8'b00011000; //    **
         11'h7d5: return 8'b00011000; //    **
         11'h7d6: return 8'b00001110; //     ***
         11'h7d7: return 8'b00011000; //    **
         11'h7d8: return 8'b00011000; //    **
         11'h7d9: return 8'b00011000; //    **
         11'h7da: return 8'b00011000; //    **
         11'h7db: return 8'b01110000; //  ***
         11'h7dc: return 8'b00000000; //
         11'h7dd: return 8'b00000000; //
         11'h7de: return 8'b00000000; //
         11'h7df: return 8'b00000000; //
         //code x7e
         11'h7e0: return 8'b00000000; //
         11'h7e1: return 8'b00000000; //
         11'h7e2: return 8'b01110110; //  *** **
         11'h7e3: return 8'b11011100; // ** ***
         11'h7e4: return 8'b00000000; //
         11'h7e5: return 8'b00000000; //
         11'h7e6: return 8'b00000000; //
         11'h7e7: return 8'b00000000; //
         11'h7e8: return 8'b00000000; //
         11'h7e9: return 8'b00000000; //
         11'h7ea: return 8'b00000000; //
         11'h7eb: return 8'b00000000; //
         11'h7ec: return 8'b00000000; //
         11'h7ed: return 8'b00000000; //
         11'h7ee: return 8'b00000000; //
         11'h7ef: return 8'b00000000; //
         //code x7f
         11'h7f0: return 8'b00000000; //
         11'h7f1: return 8'b00000000; //
         11'h7f2: return 8'b00000000; //
         11'h7f3: return 8'b00000000; //
         11'h7f4: return 8'b00010000; //    *
         11'h7f5: return 8'b00111000; //   ***
         11'h7f6: return 8'b01101100; //  ** **
         11'h7f7: return 8'b11000110; // **   **
         11'h7f8: return 8'b11000110; // **   **
         11'h7f9: return 8'b11000110; // **   **
         11'h7fa: return 8'b11111110; // *******
         11'h7fb: return 8'b00000000; //
         11'h7fc: return 8'b00000000; //
         11'h7fd: return 8'b00000000; //
         11'h7fe: return 8'b00000000; //
         11'h7ff: return 8'b00000000; //
    endcase
  endfunction

endpackage